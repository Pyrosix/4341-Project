`timescale 1ns/1ns
`include "../32_bit_or.v"

module OR_tb;
reg [31:0] a, b;
wire [31:0] s;

OR_32b test(.a(a), .b(b), .s(s));
initial begin
$dumpfile("OR.vcd");
$dumpvars(0, OR_tb);
$display("    a                               |                 b                  |  y");
$display("------------------------------------+------------------------------------+---");
$monitor("a = %b b = %b y = %b", a, b, s); 

// <# of bits>'b<binary value>
a = 32'b11111111111111111111111111111111; b = 32'b11111111111111111111111111111111; #20;  // case: both input's == 1 -> 1
a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000000; #20;  // case: both input's == 0 -> 1
a = 32'b00000000000000000000100000001000; b = 32'b00000000000000000000100000001000; #20;  // 2056 OR 2056 -> 2056
a = 32'b11111111100110001001011001111111; b = 32'b11111111100110001001011001111111; #20;  // 2147483647 == 2147483647 ? -> 1
a = 32'b11111111111111110000000000000000; b = 32'b00000000000000001111111111111111; #20;  //  [31:16] => 1's OR [15:0] 1's ? -> all 1's
a = 32'b11111111111111111111111111111111; b = 32'b00000000000000000000000000000000; #20;  //  all 1's OR all 0's -> all 1's
a = 32'b00000000000000000000000000000001; b = 32'b00000000000000000000000000000001; #20;  // 1 OR 1 ? -> 1
a = 32'b00000000000000000000000000000001; b = 32'b00000000000000000000000000000010; #20;  // 1 OR 2 ? -> 3

end
endmodule

